`ifndef DEFINES_SV
`define DEFINES_SV

//`define USE_CARRY_LOOK_AHEAD
`define ADD_SUB_OPERATOR
`define USE_DSP

`endif

